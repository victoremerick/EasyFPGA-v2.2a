/*******************************************************************
**���ǵ�FPGA������
**��վ��www.OurFPGA.com
**�Ա���OurFPGA.taobao.com
**����: OurFPGA@gmail.com���������Ƶ�̳̼�����
*****************�ļ���Ϣ********************************************
**�������ڣ�   2011.06.01
**�汾�ţ�     version 1.0
**����������   ���� 
********************************************************************/

module my_and(a,b,c);  //;������©��
input a,b;  //����a�ɿ���KEY1������0�����£�1��δ����
                   //����b�ɿ���KEY2������0�����£�1��δ����
output c;  //���c��LED��ʾ�� 0��������1��Ϩ��
assign c=a&b; //��ֱ�Ӹ�ֵ���
endmodule
